library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

use work.tipos.ALL;

entity FSM_aggregator is
        port ( 
                clk, rst                : in std_logic;

                aggregation_start       : in std_logic;

                window_done             : in std_logic;
                segment_done            : in std_logic;
                elements_done           : in std_logic;
                log_done                : in std_logic;
                padd_done               : in std_logic;

                addr_A_read_out         : out address_A;
                addr_B_read_out         : out address_B;

                data_A_select           : out padd_op_A; 
                data_B_select           : out padd_op_B; 

                k_next                  : out std_logic;
                u_next                  : out std_logic;
                m_next                  : out std_logic;
                log_next                : out std_logic;

                -- Tiene los 4 bits de control. Los 3 menos signif corresponden a las escrituras en cada componente de memoria. 
                -- El mas significativo es un data valid.
                padd_status_out         : out padd_status;
                aggregation_done        : out std_logic
);
end FSM_aggregator;

architecture Structural of FSM_aggregator is

        type states_loop is (idle, read_gs_km, read_seg_bucket, change_segment, change_element, change_to_acc, read_skskm, read_gkgkm, change_segment_b, read_skmb, read_sklog, read_wait, read_gs, wait_for_padd, endState);
        signal state_next, state_reg : states_loop;

begin

        process(clk, rst)
        begin
                if (rst = '1') then
                        state_reg <= idle;
                elsif (clk'event and clk='1') then
                        state_reg <= state_next;
                end if;
        end process;
        
        process(state_reg, window_done, segment_done, elements_done, aggregation_start, log_done, padd_done)
        begin
                state_next <= state_reg;

                case state_reg is
                        when idle =>
                                state_next <= read_gs_km when aggregation_start = '1' else
                                              idle;
                        when read_gs_km =>
                                state_next <= read_seg_bucket when window_done = '1' else
                                              read_gs_km;
                        when read_seg_bucket =>
                                state_next <= change_segment when window_done = '1' else
                                              read_seg_bucket;
                        when change_segment =>
                                state_next <= change_element when segment_done = '1' else
                                              read_gs_km;
                        when change_element =>
                                state_next <= change_to_acc when elements_done = '1' else
                                              read_gs_km;
                        when change_to_acc =>
                                state_next <= read_skskm;
                        when read_skskm => 
                                state_next <= read_gkgkm when window_done = '1' else
                                              -- Me falta un OR en esta parte (?)
                                              read_skskm;
                        when read_gkgkm =>
                                state_next <= change_segment_b when window_done = '1' else
                                              read_gkgkm;
                        when change_segment_b =>
                                state_next <= read_sklog when segment_done = '1' else
                                              read_skmb;
                        when read_skmb =>
                                state_next <= read_skskm when window_done = '1' else
                                              read_skmb;
                        when read_sklog =>
                                state_next <= read_wait when window_done = '1' else
                                              read_gs when log_done = '1' else
                                              read_sklog;
                        when read_wait =>
                                state_next <= read_sklog when padd_done = '1' else
                                              read_wait;
                        when read_gs    => 
                                state_next <= wait_for_padd when window_done = '1' else
                                              read_gs;
                        when wait_for_padd =>
                                state_next <= endState when padd_done = '1' else
                                              wait_for_padd;
                        when endState   =>
                                state_next <= state_reg;

                end case;
        end process;


        process(state_reg, window_done)
        begin

                m_next          <= '0';
                u_next          <= '0';
                k_next          <= '0';
                log_next        <= '0';

                -- Tiro valores random para inicializar esto.;
                addr_A_read_out <= g_k;
                addr_B_read_out <= bucket;
                padd_status_out <= ('0','0','0','0');

                data_A_select     <= bucket_op; 
                data_B_select     <= bucket_op;
                aggregation_done   <= '0';

                case state_reg is
                        when idle =>
                        when read_gs_km =>
                                addr_A_read_out <= g_km;
                                addr_B_read_out <= s_km;

                                data_A_select <= aux_op;
                                data_B_select <= segment_op;

                                k_next <= '1';
                                -- Escribo en aux
                                padd_status_out <= ('1','0','0','1');

                        when read_seg_bucket =>
                                addr_A_read_out <= s_km;
                                addr_B_read_out <= bucket;

                                data_A_select <= segment_op;
                                data_B_select <= bucket_op;

                                k_next <= '1';
                                -- Escribo en aux y segmento
                                padd_status_out <= ('1','0','1','1');

                        when change_segment =>
                                m_next <= '1';
                        when change_element =>
                                u_next <= '1';
                        when change_to_acc =>
                        when read_skskm =>
                                addr_A_read_out <= s_k;
                                addr_B_read_out <= s_km;

                                data_A_select <= segment_op;
                                data_B_select <= aux_op;

                                k_next <= '1';
                                -- Escribo en bucket y segmento
                                padd_status_out <= ('1','1','1','0');

                        when read_gkgkm => 
                                addr_A_read_out <= g_k;
                                addr_B_read_out <= g_km;

                                data_A_select <= bucket_op;
                                data_B_select <= aux_op;

                                k_next <= '1';
                                -- Escribo en bucket (Y aux??)
                                padd_status_out <= ('1','1','0','1');

                        when change_segment_b =>
                                m_next <= '1';
                        when read_skmb =>
                                addr_A_read_out <= s_km;
                                addr_B_read_out <= s_km_b;

                                data_A_select <= segment_op;
                                data_B_select <= aux_op;

                                k_next <= '1';
                                -- Escribo en aux y segmento
                                padd_status_out <= ('1','0','1','0');

                        when read_sklog =>
                                addr_A_read_out <= s_k;
                                addr_B_read_out <= s_k;

                                data_A_select <= segment_op;
                                data_B_select <= segment_op;

                                k_next <= '1';
                                -- Escribo en bucket y segmento
                                padd_status_out <= ('1','1','1','0');
                                if window_done = '1' then
                                        log_next <=  '1';
                                else
                                        log_next <=  '0';
                                end if;

                        when read_wait =>
                        when read_gs =>
                                addr_A_read_out <= g_k;
                                addr_B_read_out <= s_k;

                                data_A_select <= bucket_op;
                                data_B_select <= segment_op;

                                k_next <= '1';
                                -- Escribo en bucket
                                padd_status_out <= ('1','1','0','0');

                        when wait_for_padd =>
                        when endState =>
                                aggregation_done <= '1';
                end case;
        end process;

end Structural;
